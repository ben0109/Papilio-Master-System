library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library UNISIM;
use UNISIM.vcomponents.all;

entity vdp_vram is
	Port (clk		: in  STD_LOGIC;
		cpu_WE		: in  STD_LOGIC;
			cpu_A		: in  STD_LOGIC_VECTOR (13 downto 0);
			cpu_D_in	: in  STD_LOGIC_VECTOR (7 downto 0);
			cpu_D_out: out STD_LOGIC_VECTOR (7 downto 0);
			vdp_A		: in  STD_LOGIC_VECTOR (13 downto 0);
			vdp_D_out: out STD_LOGIC_VECTOR (7 downto 0));
end vdp_vram;

architecture Behavioral of vdp_vram is
begin
	RAMB16_S1_inst0 : RAMB16_S1_S1
	generic map (
		INIT_00 => X"0000000000000000000000000070000000000000000000000000070007006000",
		INIT_01 => X"00700000577750770000007000000000700055ee000007000000770077000000",
		INIT_02 => X"0000000000000000000000000070000000000000000000000000070007000000",
		INIT_03 => X"007000000677b07700000070000000000007bb33000007000000770077000000",
		INIT_04 => X"0000000000000000000007000070000000000000000000000000007007000000",
		INIT_05 => X"0000000000000000007000000000070000000000000000000000700000070000",
		INIT_06 => X"0000000066666600066600066666666600000000000000007000000000000007",
		INIT_07 => X"06666666eeeeeee0666666666066666606666666606666776600066666777600",
		INIT_08 => X"0000000000000000555555555777775530000000eeee0333eee0333366667760",
		INIT_09 => X"666666666666666600666666666777760000000000000000bbbbbbbbb77777bb",
		INIT_0A => X"eee06666e0eee06633330eee33333333eeeeeeee0000eee066666000eeeeeeee",
		INIT_0B => X"066666660666666666666666e0066666066666660000066666666000eee00000",
		INIT_0C => X"eeeeeeee333330000000000030eeeeeeeeeeeeeeeeeee000000e06666776000e",
		INIT_0D => X"66000000666666000000eeee60eeeeee6000eeeeeeeee06666600eee60eeeeee",
		INIT_0E => X"3330000000000000ee003333eeeeeeeee000000006666666eee00666eeeeeeee",
		INIT_0F => X"666666766666666600066677666666606006666666666666eeeeeeee03333333",
		INIT_10 => X"00000000eee03330eeeeeeee66000eee666000ee006666007606666666000006",
		INIT_11 => X"6666606666666066e066666666600006e060000666666666eeeeeeee33333333",
		INIT_12 => X"00000000303330eeeeeeeeee0eeee66600000666e00000006666667766006666",
		INIT_13 => X"66666606eeeeeeeee00006666666600006666666eeeeeeee330e000e00000033",
		INIT_14 => X"000003330033330eeeee000000666666eeeeeeee66606666ee06666666666666",
		INIT_15 => X"0eee066630ee0666eeeeeeee33333306eeeeeeee33333300eeeeee0300000000",
		INIT_16 => X"0000000000000000eeeeee0e6666000e666660006660000e66666666eeeeeeee",
		INIT_17 => X"0000333300003333000033300003330e000000033330eeee00030033003330ee",
		INIT_18 => X"00003333000000003330eeeeeeeeee060eeee066eeee066600eeee06033330ee",
		INIT_19 => X"666666600000666000006660eeeeeeee00000003033330ee00333333033330ee",
		INIT_1A => X"0000000000000000666666606666666000006660000066606666666000000000",
		INIT_1B => X"0000000066666666666666660000000060000000666666666666666060666666",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"00000000eee03333000000333330000000000000067000660000000000000000",
		INIT_1E => X"00000000000000000000000000000000eeeeeeeeee000000eee0000000000000",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0000000000000000000000000000000000000000000400000000000000000000",
		INIT_21 => X"0000000000000000003020000000000000000000000000000000000000000000",
		INIT_22 => X"0000001000000004000000000000000000000000000000000000000000030000",
		INIT_23 => X"0000000000000000400000040000000000000000000000000000000000000000",
		INIT_24 => X"0000000000000000000000020000000030000000020200000000000000000200",
		INIT_25 => X"0000000000040000000000000001040000000000000000000000000000000000",
		INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => X"0030000000020000000000000002000000000000000000000000000000000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000000009000090000000000009009000090900000000000000000000000000",
		INIT_2D => X"0000000000000000000000000000000000009000009000900000000000000000",
		INIT_2E => X"0000009900990000009990000009000000990009090009900900000000099900",
		INIT_2F => X"0000099099999999000000000000000000000000000000000009999000990000",
		INIT_30 => X"0999900900000009090090090009990000900090009909900999990000999900",
		INIT_31 => X"0099999009999999099999990900000009000009009999990900000909999999",
		INIT_32 => X"0999999900009999009999990000000900990000090099900909999000009990",
		INIT_33 => X"0000000000000000000000000000000000000000090000990000099909900099",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"5555555500000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"febfebebebbfebfebafeebfbbbefaeffabfaeeefebebbeafaaabebbfeaaebfaa",
		INIT_39 => X"abefeefbbfffffefbafaebfaaeaeefbebebabaffabffaebbefafbbbebbbeeaab",
		INIT_3A => X"abeafaabbfbffeabefabaabffaafbfaafebeafaeeaaaabfafffebeeabffbeaff",
		INIT_3B => X"febabbaeeaaaaabaefafbeaffbfbbaebebefeffbaeeafbeebafeffeaaeeeeffe",
		INIT_3C => X"febfaffeeaeaabfebafeffeaaffaeaffabebfafbbffffeafaaabebbfeaaebfaa",
		INIT_3D => X"abefeefbbfffffefbafaebfaaeaeefbebebabaaefbbfaebbefabaabffbbbbaab",
		INIT_3E => X"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
		INIT_3F => X"0550005000000055005500000000000000000000000000000ffc3f3fff0f00ff"
	)
	port map (
		CLKA => clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(0 downto 0),
		DOA => cpu_D_out(0 downto 0),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(0 downto 0),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst1 : RAMB16_S1_S1
	generic map (
		INIT_00 => X"0000000000000000000000000007000000000000000000000000700700066600",
		INIT_01 => X"0070000067775077000000077000000077775500000007000000000700000000",
		INIT_02 => X"0000000000000000000000000007000000000000000000000000700700006600",
		INIT_03 => X"007000000667b07700000007700000007777bb00000007000000000700000000",
		INIT_04 => X"0000000000000000000007000070000000000000000000000000000770000000",
		INIT_05 => X"0000000000000000007000000770070000000000000000000000700007070000",
		INIT_06 => X"6666660066677760666666666666666600000077770000007000000000777007",
		INIT_07 => X"66666666eeee000066666600606666666666666666066777606666666666760e",
		INIT_08 => X"000000ffff000000555555555777775533300000eeeee033eee0000066666760",
		INIT_09 => X"00006666666666666606666066666677000000aaaa000000bbbbbbbbb77777bb",
		INIT_0A => X"eee06666030eee000333300e33333333eeeeeeee00000ee066666666eeeeeeee",
		INIT_0B => X"066660006666666606666666e0666666e06666660066666666666000eeeeee00",
		INIT_0C => X"eeeeeeee300000000000033330eeeeeeeeeeeeee0eee00006000e06666666000",
		INIT_0D => X"776600006666660e6000eeee0eeeeeee6000eee0eeeee06666600eee0eeeeeee",
		INIT_0E => X"3300000000000000eeee0333eeeeeeee00000000e0666666eee006660eeeeeee",
		INIT_0F => X"66666666666666600ee066676666600000e0666666666660eeeeeeee03333333",
		INIT_10 => X"00000000eee03330eeeeeeee766000ee666000ee667777607760666760666666",
		INIT_11 => X"6666606666660666e0666660666660000666666666666666eeeeeeee33333333",
		INIT_12 => X"00000000003330eeeeeeeeee00ee066760006666000000066666666666660666",
		INIT_13 => X"66666660eeeeeeee0006666666666000e00666660eeeeeee3300330e00000003",
		INIT_14 => X"000033330033330eeee0000006666666eeeee00066006666ee00000066666666",
		INIT_15 => X"eeee06663300e066eeeeeeee33000006eeeeeeee33333333eeee003300000000",
		INIT_16 => X"0000000033300000eeeeeeee67766000666666006660000e66666666eeeeeeee",
		INIT_17 => X"00033330000003330000333000033330000003333330eeee0000333300033300",
		INIT_18 => X"0000033300000333330eeeeeeeeee06630eee066eeeee066330000000333330e",
		INIT_19 => X"666660600000666000006660eeeeeeee00000003333330ee0003333303330eee",
		INIT_1A => X"6000000000000000006666606666660000006660000066606666666066000000",
		INIT_1B => X"0000000066666000066666660000000000000000666666666666666666666666",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"00000000eeee0333000033300300000000000000066000660000000000000000",
		INIT_1E => X"00000000000000000000000000000000eeeeeeeee00660000000000000000000",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0000000400000000000000000000000000000000000000000000000000000000",
		INIT_21 => X"0000310000000000400000000101000000000000020000000000200000010000",
		INIT_22 => X"0000000000000000003000000001000000000000000000000000000000000000",
		INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_24 => X"0000000000002000000000000000000020100000000000000040000000000000",
		INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => X"0000000000000000000030000001000000000000000400000000000000000000",
		INIT_27 => X"0000000000000000000000000000000000000004000000000000000000000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000000009900990000000000090909009999999000009990000099000000000",
		INIT_2D => X"0000000000000000000090000000000000009000009909900000000000000000",
		INIT_2E => X"0000099909999009099999090999999909999099090099990900000000999990",
		INIT_2F => X"0000999999999999000909000000000000000000000000000099999909990990",
		INIT_30 => X"0999900900009009090090090099999009900099099999990999999009000090",
		INIT_31 => X"0999999909999999099999990900000009900099099999990900000909999999",
		INIT_32 => X"0999999900099999099999990000000909999090099099990099999900099999",
		INIT_33 => X"9900000000090000000000000000000000009000090009990000999909990999",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"5555555500000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"5150401450041500015400051104111514414511110015410001400014441051",
		INIT_39 => X"5015151040540045541504045400140140414014015540105551415050440004",
		INIT_3A => X"0545441515415454111010110555014015140505114511440000011554400551",
		INIT_3B => X"5150514155015500444545545004511554515054041044011055544010045005",
		INIT_3C => X"0405141400540055541110045550144041000001514510145554155541114504",
		INIT_3D => X"0540404515015510014051510155415415141505005015450001010014401551",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"d88d88d8dd8888d888dd888d8888dddd0000000000000000ffc00ff0ffcfffff"
	)
	port map (
		CLKA => clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(1 downto 1),
		DOA => cpu_D_out(1 downto 1),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(1 downto 1),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst2 : RAMB16_S1_S1
	generic map (
		INIT_00 => X"0000000000000000e0000000000700000000000000000000000070700006660e",
		INIT_01 => X"0070000066775057000000000777000077755000007007000000777000000000",
		INIT_02 => X"0000000000000000000000000007000000000000000000000000707006066033",
		INIT_03 => X"00700000066bb0b70000000007770000777bb000007007000000777000000000",
		INIT_04 => X"0000000000000000000000777700000000000000000000000000000000000000",
		INIT_05 => X"0000000000000000000700000000700000000000000000000000070000700000",
		INIT_06 => X"6666666066667776666666666666666600007700007700000700000007770070",
		INIT_07 => X"666666660000000066600000606666666666666666066666066666666666660e",
		INIT_08 => X"0000ff5555550000055555555777775033333000eeeee033eeeeeeee06666666",
		INIT_09 => X"000000660066666666600006666666660000aabbbbbb00000bbbbbbbb77777b0",
		INIT_0A => X"eee066663330eeee0333333033333333eeeeeeee66000eee66666666eeeeeeee",
		INIT_0B => X"e0600000666666660666666600666666e06666666666666666666660eeeeee06",
		INIT_0C => X"eeeeeee000000000000333330eeeeeeeeeeeeeee0eee06666000006666666000",
		INIT_0D => X"677660006666660e6000eeeeeeeeeeee6000eee000eee06666600eeeeeeeeeee",
		INIT_0E => X"3000000000000000eeeee033eeeeeeee06666600e0666666eeeee0660eeeeeee",
		INIT_0F => X"006666660000000e0ee0666600000000000006660000000eeeeeeeee03330000",
		INIT_10 => X"00000000ee03330eeeeeeeee776000ee66600eee666667766660666600000666",
		INIT_11 => X"6666066600006666e0666660667776600666666000000000eeeeeeee33333333",
		INIT_12 => X"00000000ee03330eeeeeeeee00ee066666666666000066666666666600666000",
		INIT_13 => X"66666666eeeeeeee0666666666666000eee0000030eeeeee3033330e00000000",
		INIT_14 => X"000333300003330eee06666066666666ee000000000666660000000066660000",
		INIT_15 => X"eeee066633330066eeeeeeee00eeee06eeeeeeee000033330000333333300000",
		INIT_16 => X"0000000333333000eeeeeeee66776000000006666666000e666666660eeeeeee",
		INIT_17 => X"00033330000000330000330e00003330000333303330eeee0003333300033333",
		INIT_18 => X"0000003300033333330eeeeeeeeee06630eee000eeeee0663333330000333330",
		INIT_19 => X"660000006666666000006660eeeeeeee00000003333330ee0000033303330eee",
		INIT_1A => X"6666666600000000000666606666660000006660000066606666666066666060",
		INIT_1B => X"0000000066660000066666666000000000000000666666666666666666666666",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"00006666eeee0333770333307000000000700000666666660000000000000000",
		INIT_1E => X"00000000000000000000000000000000eeeeeeeee00666663006666700006677",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0000000000000000000000030000003000300000000000000000000000000000",
		INIT_21 => X"0000000000002000000000000000300000000000000000000000000000040000",
		INIT_22 => X"0000000000000000000000000000000000000000030000000000000000000000",
		INIT_23 => X"0000000000000000400000000402000000000000000000000000020000000000",
		INIT_24 => X"4000000000000000000000000000000000000000000000000010000000000000",
		INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => X"0000000000000000000000000000000000000000000000000000000000004000",
		INIT_27 => X"0000000000000000000000000000000000000000000000000000040000000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000000000999900000000000999999909999999000009990000999900000000",
		INIT_2D => X"0000000000000000000090000990000000999990000999000000000000000000",
		INIT_2E => X"0000990909009009090009090999999909009999090999090999999909000999",
		INIT_2F => X"0909909999999999000909000000000009900990099009900990900909099009",
		INIT_30 => X"0900900900009009090090090990009909000009090090090009009990000009",
		INIT_31 => X"0900000900999000000099900900000009990990090000000999999900009000",
		INIT_32 => X"0099900000999000090000000999999909009099099990090999000900090009",
		INIT_33 => X"9900990000999000000090000000900000009000090099990999900000999990",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"5555555500000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"0555505140104401410550014010514551414511400455145551501554414455",
		INIT_39 => X"1441550105551555040051541544055400514501455001151110145451404540",
		INIT_3A => X"0010041501455054141150540500150504545101115101400005454001100100",
		INIT_3B => X"4111044450544045414504014411540155041040045054500141001110054015",
		INIT_3C => X"5405114141115101404405105050415045150150440455555550101540055404",
		INIT_3D => X"4454401145011510501555504144115540100545550541054440010445545544",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"a5a505a0f505a0f005a5f000f5f5f5f5000000000000000033c33c3fcfccffff"
	)
	port map (
		CLKA => clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(2 downto 2),
		DOA => cpu_D_out(2 downto 2),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(2 downto 2),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst3 : RAMB16_S1_S1
	generic map (
		INIT_00 => X"0000000000000000e550000000007000000000000000000000070070005550ee",
		INIT_01 => X"00070000666750ee0000000000007777e5555000077070007777000000000000",
		INIT_02 => X"0000000000000000bbb0000000007000000000000000000000070070666bb033",
		INIT_03 => X"00070000066b66330000000000007777bbbbb000077070007777000000000000",
		INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_05 => X"0000007777000000000077000077000000000000000000000000007777000000",
		INIT_06 => X"6666666066666676666666606666666600770000000077000700000000000070",
		INIT_07 => X"66666660000000660000000006600666666666666606666600000666666660ee",
		INIT_08 => X"00ff555555555500055555555577755033333300eeeee033ee00000e06666666",
		INIT_09 => X"000000060e066666666666666666666600aabbbbbbbbbb000bbbbbbbbb777bb0",
		INIT_0A => X"eee06666330eeeee0033333330000033eeeeeeee766000ee666666660eeee000",
		INIT_0B => X"e000000066666660e066666606666666e06666666666666666666666eeeee066",
		INIT_0C => X"eeeeee0300000000003333330eeeeeeeeeeeeeee00e066670000066666666600",
		INIT_0D => X"66666000666660ee6600eeeeeeeeeeee6000ee06000eee0666600eeeeeeeeeee",
		INIT_0E => X"0000000000000000eeeeee03eeeeeeee66677660e0666666eeeee0660eeeeeee",
		INIT_0F => X"0e0666660000000e00e066660666660000000666eeeeeeeeeeeeeeee03330000",
		INIT_10 => X"333000000033330eeeeeeee0676000ee66600eee666666666660666600000000",
		INIT_11 => X"0000666066666600e06666606667776606666660eeeeeeeeeeeeeeee00333330",
		INIT_12 => X"00000033ee033330eeeeeeee000e066666666666600000066600066600000000",
		INIT_13 => X"66666666eeeeeeee6666666666666000eeeeeeee330eeeee0333330e00000000",
		INIT_14 => X"0003330e00033330e06677666666666600000006ee0666660000000066600ee0",
		INIT_15 => X"eeee0666333330060eeeeee0eeeeee06eeeeeeeeeeee00333333333333330000",
		INIT_16 => X"0000003300333330eeeeeeee666760000000006666660000666600003000eee0",
		INIT_17 => X"00033330000000000003330e000033330033330e3330eeee0003330000003333",
		INIT_18 => X"0000000000333300330eeeeeeeeee06630eee000eeeee0663333330000033333",
		INIT_19 => X"000000006666666000066660eeeeeeee00000003333330ee0000333303330eee",
		INIT_1A => X"6666666600000000000066606666600066666660000066606666666066666660",
		INIT_1B => X"0000000066600000006666666666666600000000666666666066666666666660",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"00066666eeee0333667033306700000006670000666666660000000000000000",
		INIT_1E => X"00000000000000000000000000000000eeeeeeeee00066663006666600066666",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0000000000000000000000000040000000000000000000000000000000000000",
		INIT_21 => X"0002000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => X"0000000000000000000000000000000000000000001000000003000000000000",
		INIT_23 => X"0400000000200000000000010000000000000000000000000000000400000000",
		INIT_24 => X"0000000000000000010000000000000000000000000000000000000000000000",
		INIT_25 => X"0000000000002000000000000000000000000000000000000000000010000000",
		INIT_26 => X"0000000000000000000000000000000000000000001000000000000000000000",
		INIT_27 => X"0400000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000009900099000000000000090909000090900000000000000999900000000",
		INIT_2D => X"0000000000000000000090009990000000999990099999990000000000000000",
		INIT_2E => X"0999900909009009090009090009009909009909090990090999999909000009",
		INIT_2F => X"0909009999999999000909000000000099900990099009900900900909099009",
		INIT_30 => X"0900000900009009090090090900000909000009090090090009000990900909",
		INIT_31 => X"0900000900099900000999000900000000999900090000000999999900009000",
		INIT_32 => X"0009990009990000090000000999999909009009009900090909000900090009",
		INIT_33 => X"0000990009999900000990000000990000009000090999090999900000099900",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"5555555500000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"1015411050045540500010110040105104404154004145054044444004105010",
		INIT_39 => X"0511514450554110411044540444504401505510414445115450005410001015",
		INIT_3A => X"0104545444511405550451400050444011414105501051545151501114114001",
		INIT_3B => X"5510401111441001114451445544115445455450510500404505450501111511",
		INIT_3C => X"4410540515500415045145514111150141515044050514501510511545050514",
		INIT_3D => X"4045111105541400104511054511011154444044111110541014551055501140",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"4ee4411be4444ee4444eb441ee44bb1100000000000000000ff00fc0cf0cffff"
	)
	port map (
		CLKA => clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(3 downto 3),
		DOA => cpu_D_out(3 downto 3),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(3 downto 3),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst4 : RAMB16_S1_S1
	generic map (
		INIT_00 => X"7777000000000000777550000000700000000000000077770007000006555057",
		INIT_01 => X"000700006665550e0000000000000000e5500000070070000000000000000000",
		INIT_02 => X"7777000000000000777bb000000070000000000000007777000700006667b0b7",
		INIT_03 => X"0007000006b666000000000000000000bbb00000070070000000000000000000",
		INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_05 => X"0000770000770000000000777700000000000077770000000000000000000000",
		INIT_06 => X"0000006066666666666666000000066607000000000000700077000000007700",
		INIT_07 => X"6660000e0006666600000000660ee06666660000606666660000006600000eee",
		INIT_08 => X"0f55555555555550005555555555550003333330eeeee033e000000006666666",
		INIT_09 => X"666600000060000066666666660066660abbbbbbbbbbbbb000bbbbbbbbbbbb00",
		INIT_0A => X"eee06666330eeeee000333330eeeee00eeeeeeee776000ee666666660e000000",
		INIT_0B => X"e000066666666660e066666606666666ee0666666666666666666666eeeee066",
		INIT_0C => X"eeee00330000000003333300eeeeeeeeeeeeeeee00e066660000066666666600",
		INIT_0D => X"6666660000000eee6600eeee0eeeeeee600eee060000ee0666600eeeeeeeeeee",
		INIT_0E => X"0000000000000000eeeeeee0eeeeeeee66667760ee066600eeeeee06eeeeeeee",
		INIT_0F => X"0006666666660000000066660666666600006666eeeeeeeeeeeeeeee33330000",
		INIT_10 => X"33333033333330eeeeeeeee0666000ee6660eeee066666606006666600000000",
		INIT_11 => X"6666666066000006e06666606666677606666660eeeeeeeeeeeeeee000000000",
		INIT_12 => X"00003333eee03333eeeeeeee000e066666666666000000006000e06660000000",
		INIT_13 => X"66666666eeeeeeee6666666666666600eeeeeeee330eeeee0000033000000000",
		INIT_14 => X"003330ee03333330e06667766666666600066660ee0666660666666666600ee0",
		INIT_15 => X"eeee066633300ee030eeeee0eeeeee06eeeeeeeeeeeeee033333330033330000",
		INIT_16 => X"00000033ee003333eeeeeeee6666600066000066666600000000eeee33330000",
		INIT_17 => X"00033330000000030003330e00000333033330ee33330eee003330ee00000033",
		INIT_18 => X"00000000033330ee330eeeeeeeeee0660eeee066eeeee0660003330e00000333",
		INIT_19 => X"000000006666666000000000eeeeeeee00000333333330ee00033333033330ee",
		INIT_1A => X"6666666666600000000066606660000066666660000666600000006066666660",
		INIT_1B => X"0000666666600000000066666666666600000000600000000066000666660000",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"0000666600000033066033006660000000600000666666600000000000000000",
		INIT_1E => X"00000000000000000000000000000000ee000000e00660660000000000006666",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0000000000000000000000000000000000010003000000000000000000000000",
		INIT_21 => X"0000000000300000000000000000000000000000000020000003000000000000",
		INIT_22 => X"0001000000000000010000000000000000000000000040200000000000000020",
		INIT_23 => X"0000000000000000000000000000000000000000000000000004000000000000",
		INIT_24 => X"0000000000000030000000000000103000000000000000000000000000000000",
		INIT_25 => X"0000000000000002000000000000000000000000100000200000000000000000",
		INIT_26 => X"0000000000000000000000000000000000000000000000000000003000000001",
		INIT_27 => X"0000000000000002000000000000000000000000000000000000000000000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000099900999900000000000999999909999999000009990990999000000000",
		INIT_2D => X"0000000009900000000090009000000000009000099999990000000000000000",
		INIT_2E => X"0999000909009099090009090009099009009009099990090900009009900009",
		INIT_2F => X"0909009999999999000909000000000090000000000000000900900909009909",
		INIT_30 => X"0990009900009009090090090900000909900099090090090009009990900909",
		INIT_31 => X"0900000900009990000099900900000000099000090000000900000900009000",
		INIT_32 => X"0099900000999000090000000000000909009009000900090900000900090009",
		INIT_33 => X"0000000000090000009999900999999000999990099990090000999900999990",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"5555555500000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"5455bbafaaaa8400047baabefabeea45102aaaaaabaeba514014155544501511",
		INIT_39 => X"40101140554554511001105114111005005100abaaa44504444befaaaaeaad50",
		INIT_3A => X"5050041141005110144010140444044004101054110145045400014150441115",
		INIT_3B => X"1405145441404155044104554005041150511540054050414041150040051544",
		INIT_3C => X"0144101555155504111410005050105440040501110154104415155114440104",
		INIT_3D => X"1145004041545140115510414411000545441140115444515554011510500101",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"500f04145f05505a05054f04ffaa1144000000000000000030cc3ccff3cf3cc3"
	)
	port map (
		CLKA => clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(4 downto 4),
		DOA => cpu_D_out(4 downto 4),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(4 downto 4),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst5 : RAMB16_S1_S1
	generic map (
		INIT_00 => X"0000777000000000777750000000070000000000077700000070000006655077",
		INIT_01 => X"0000700006066055000000000000000000000000000700000000000000000000",
		INIT_02 => X"00007770000000007777b000000007000000000007770000007000006677b077",
		INIT_03 => X"0000700000b666bb0000000000000000b0000000000700000000000000000000",
		INIT_04 => X"0000007777000000000000000000000000000000000000000000000000000000",
		INIT_05 => X"0007000000007000000000000000000000000700007000000000000000000000",
		INIT_06 => X"000000000066666666666600eeeee00007000000000000700000770000770000",
		INIT_07 => X"000eeeee666666660666666660000066000000000666006600000006eeeeeeee",
		INIT_08 => X"0f555555555555500000555555550000e0033330eeee033300000000e0666666",
		INIT_09 => X"677766000066666666666666600e00000abbbbbbbbbbbbb00000bbbbbbbb0000",
		INIT_0A => X"eee06666330eeeee00000333eeeeeeeeeeeeeeee6760000e6666666000000000",
		INIT_0B => X"e006666666666660ee06666606666666ee0660006666666666666666eeee0666",
		INIT_0C => X"ee00333300000000333300eeeeeeeeeeeeeeeeee00e066660000006666666660",
		INIT_0D => X"6666660000eeeeee6600eeee00eeeeee600ee06660000ee06660eeeeeeeeeeee",
		INIT_0E => X"0000000033300000eeeeeeeeeeeeeeee66666760ee066000eeeeee06000eeeee",
		INIT_0F => X"0066666666666600000666660666677666666666eeeeeeeeeeeeeeee33330000",
		INIT_10 => X"0033330333300eeeeeeeeee0666000ee6600eeee000060000666600666666000",
		INIT_11 => X"6666660000000666e06666666666666660666606eeeeeeeeeeeeeee000000000",
		INIT_12 => X"00033330eeee0033eeeeeeee000e066666666666000000006000060076600066",
		INIT_13 => X"00666660eeeeeeee6666666666666666eeeeeeee330eeeee0000033000000000",
		INIT_14 => X"003330ee33330000e06666766666666666666000ee0666666666667766600e06",
		INIT_15 => X"eeee0666330eeeee3300ee06eeeeee06eeeeeeeeeeeeee030000000033330000",
		INIT_16 => X"00000033eeee0333eeeeeeee666660007660006666660006eeeeeeee3300ee06",
		INIT_17 => X"00033330000000330003330e0000003303330eee03330eee003330ee00000000",
		INIT_18 => X"0000000003330eee00eeeeeeeeeee066eeee0667eeeeee06003330ee00000033",
		INIT_19 => X"000666606666666000000000eeeeeeee000333333333330e00033330003330ee",
		INIT_1A => X"6666666666666000000066600000000066666660000000000000000000666660",
		INIT_1B => X"0066666666600000000000006666666600000000000000000066000060000000",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"0000000000000003066033006700000000000070000000000000000000000000",
		INIT_1E => X"00000000000000000000000000000000e0000000e00660660000000000000000",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0000004000000000000000000000000000000000000000000000000000000000",
		INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => X"0000000000000000000000100000000000000000000000000000000000000000",
		INIT_23 => X"0000000000000000000000000000000000000000000000000000001000000000",
		INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_25 => X"0004404000000000000000000000000004000000000000000000000000000000",
		INIT_26 => X"0000200000000000000000000000000000000000000000000000000000000000",
		INIT_27 => X"0000000000002000000000000000000000040000000000000000000000000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000090009900990000000000090909009999999000009990990000000000000",
		INIT_2D => X"0000000009900000000090000000000000009000000999000000000000000000",
		INIT_2E => X"0000009909999990099009990009990009900009099900990900000000999990",
		INIT_2F => X"0000099999999999000909000000000000000000000000000900999909009999",
		INIT_30 => X"0099999009999999099999990999999900999990099999990999999090099009",
		INIT_31 => X"0999999909999999099999990999999909999999099000000900000909999999",
		INIT_32 => X"0999999900099999099999990000000909909999099999990999999909999999",
		INIT_33 => X"0000000000090000000990000000990000099900099900090000099909990999",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"5555555500000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"1151040004401554544405400400005554041000041040445114154441544500",
		INIT_39 => X"4515055451414410101441455505444000105140100044511114000104010055",
		INIT_3A => X"0115015005055505501450500105411140504004051555045551050141155541",
		INIT_3B => X"4154100541055451041555040544501544515555551545540150101415544014",
		INIT_3C => X"1554011101544144404544154150414010115441115450514100015055544101",
		INIT_3D => X"5155004055545015044455411111405450114514554451050500004511405051",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"aaffaaeaffaffaaaafffaaaa5500110000000000000000000f3f03f000f03c00"
	)
	port map (
		CLKA => clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(5 downto 5),
		DOA => cpu_D_out(5 downto 5),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(5 downto 5),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst6 : RAMB16_S1_S1
	generic map (
		INIT_00 => X"0000000700000000700055000000070000000000700000000070000006675077",
		INIT_01 => X"0000700000006600000000000000000000000077000700000000000000000000",
		INIT_02 => X"00000007000000000007bb00000007000000000070000000007000006777b077",
		INIT_03 => X"0000700000006000000000000000000000000077000700000000000000000000",
		INIT_04 => X"0000070000700000000000000000000000000007700000000000000000000000",
		INIT_05 => X"0070000000000700000000000000000000007000000700000000000000000000",
		INIT_06 => X"00000000ee06666666666000eeeeeeee70000000000000070000007777000000",
		INIT_07 => X"eeeeeeee6666666666667777600006660000000066600e0666666000eeeeeeee",
		INIT_08 => X"f5555555555555550000005555000000eee03333eeee033006666600e0666666",
		INIT_09 => X"66677760006666666660000060006666abbbbbbbbbbbbbbb000000bbbb000000",
		INIT_0A => X"eee066663330eeee00000000eeeeeeeeeeeeeeee6666000e6660000e00000666",
		INIT_0B => X"0066666666666660ee00066606666666ee0000006666660006666666eeee0666",
		INIT_0C => X"00333333000000003330eeeeeeeeeeeeeeeeeeee000e06666660006666666660",
		INIT_0D => X"66666600000eeeee660eeeee000eeeee60eee06666000eee6600eeeeeeeeeeee",
		INIT_0E => X"0000000033333000eeeeeeeeeeeeeeee06666666ee066006eeeeeee000000eee",
		INIT_0F => X"6666666666677760666666660666667766666666eeeeeeeeeeeeeee033330000",
		INIT_10 => X"ee033303000eeeee0000eeee666000ee0000000e00000000606600e066677760",
		INIT_11 => X"66666600ee006666000066660066666666000066eeeeeeee0eeeee0300000000",
		INIT_12 => X"3303330eeeeeee00eeeeeee0000e066600000000666666606000066677660666",
		INIT_13 => X"ee00000eeeee00006666660066666666eeeeeeee330eeeee0000033300000000",
		INIT_14 => X"003330ee3000eeeee06666660000000066660006ee0666666666666666600006",
		INIT_15 => X"0eee066630eeeeee33330006eeeeee06eeeeeeeeeeeeee030000000033300000",
		INIT_16 => X"00000003eeeee033000000ee666660007760000066666666eeeeeeee30eee066",
		INIT_17 => X"00033333000003330003330e0000000333330eee033330ee003330ee00000000",
		INIT_18 => X"000000003330eeeeeeeeeeeeeeeee066eeee0666eeeeee06033330ee00000333",
		INIT_19 => X"000066606666666000000000eeeeeeee003333300333330e0033330e0033330e",
		INIT_1A => X"6666666666666600000666600006666066666660000000600000000000666660",
		INIT_1B => X"0666666666660000000000006666666660000000600000000066000000000000",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"0000000066677703066030006670000007000067000000000000000000000000",
		INIT_1E => X"00000000000000000000000000000000e0066666e00666660006666600000000",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0000300000000000000000003000000000000000000002000001000000000000",
		INIT_21 => X"0000000000000000000000000000000000010000000000000000000000400000",
		INIT_22 => X"0000000000000003000000000040000100000000000000000000000000000000",
		INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_24 => X"0000000000000003000000000000000003000000000000000000000000000000",
		INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => X"0020000000000000000000000000000000000000000000000000300000000000",
		INIT_27 => X"0000000000000000000000000000000000000000000002000000000000020000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000000009000090000000000000090000090900000000000000000000000000",
		INIT_2D => X"0000000000000000000000000000000000000000009909900000000000000000",
		INIT_2E => X"0000009900999900009009990009900000900000099000900000000000099900",
		INIT_2F => X"0000099099999999000000000000000000000000000000000000099000990990",
		INIT_30 => X"0009990009999999099999990999999900099900099999990999990009000090",
		INIT_31 => X"0099999009999999099999990999999909999999009000000000000009999999",
		INIT_32 => X"0999999900009999009999990000000000900990099999990099999009999999",
		INIT_33 => X"0000000000090000000090000000900000009000099000090000000009900099",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"5555555500000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"0000040004400000000405400400000000041000041040000000000000000000",
		INIT_39 => X"0000000000000000000000000000000000040040100010000004000104010000",
		INIT_3A => X"0000000000000000000004000000000000000000000000010000000000000000",
		INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => X"0000000000000000000000000004000000000000000000000000000000000040",
		INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"00500055000550050500550000554455000000000000000000ffcf00ffcf3cff"
	)
	port map (
		CLKA => clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(6 downto 6),
		DOA => cpu_D_out(6 downto 6),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(6 downto 6),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst7 : RAMB16_S1_S1
	generic map (
		INIT_00 => X"0000000077000000555555e00000070000000077000000000070000006775055",
		INIT_01 => X"0000070000000000000000000000000000007770007000000000000000000000",
		INIT_02 => X"0000000077000000bbbbbb3000000700000000770000000000700000b777b0bb",
		INIT_03 => X"0000070000000000000000000000000000007770007000000000000000000000",
		INIT_04 => X"0000070000700000000000000000000000000070070000000000000000000000",
		INIT_05 => X"0070000000000700000000000000000000007000000700000000000000000000",
		INIT_06 => X"66660000e060666000000666eeeeeeee70000000000000070000000000000000",
		INIT_07 => X"eeeeeeee6666666606666677006666660000666666000006777766000000000e",
		INIT_08 => X"f5555555557775550000000000000000eeee0333eeee03336667766000666666",
		INIT_09 => X"66666766006666660006666060006666abbbbbbbbb777bbb0000000000000000",
		INIT_0A => X"eeee06663330eeee00000000eeeeeeee000eeee066660000000eeeee00666666",
		INIT_0B => X"0666666666666660e000000006666666e000000066666000e0066666eeee0666",
		INIT_0C => X"3333333000000000330eeeeeeeeeeeeeeeeeee00000e06667766000066666666",
		INIT_0D => X"66666600000eeeee660eeeee0000eeee0eeee06676600eee660eeeeeeeeeeeee",
		INIT_0E => X"0000000000333303eeeeeeeeee00000e06666666eee00666eeeeeee0000000ee",
		INIT_0F => X"6666666666666776666666666666666766666666eeeeeeeee000000333300000",
		INIT_10 => X"eee03330eeeeeeee00000eee666000ee00000000600000006660000066666776",
		INIT_11 => X"66666066ee06666600000066e006666066666666eeeeeeee3000003300000000",
		INIT_12 => X"303330eeeeeeeeeeeeeeee0000000666eeee0000666677766000666667766066",
		INIT_13 => X"eeeeeeeeee0000006666600066666666eeeeeeee330eee0e0000003300000000",
		INIT_14 => X"003330ee0eeeeeee00666666eeeeeeee66600666ee0666666666666666660006",
		INIT_15 => X"0eee06660eeeeeee03333306eeeeeee0000000eeeeeeee030000000000000033",
		INIT_16 => X"00000000eeeeee000000000e66666000666000ee66666666eeeeeeee0eeee066",
		INIT_17 => X"00003333000003330003330e000000003330eeee00333300003330ee00000000",
		INIT_18 => X"000000003330eeeeeeeeeee0eeeee066eeee0666eeeeee06033330ee00003333",
		INIT_19 => X"000066600000666000000000eeeeeeee0333330e03333330003330ee00033330",
		INIT_1A => X"6000000066666600006666600000666066666660666666600000000066666660",
		INIT_1B => X"0666666666666000000000006666666666666666666600000066000600000000",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"0000000066666603300300006600000006700067000000000000000000000000",
		INIT_1E => X"00000000000000000000000000000000ee066666ee0066600006666600000000",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0030000030000000000000000000000000000000000000000000000000000000",
		INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => X"0000000000000200000000000003000003000000000000000000000010000000",
		INIT_23 => X"0000000010000300040000001000000000000000000000000000000000000000",
		INIT_24 => X"0000000000000000000000000000000000003000000000000000000000000000",
		INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => X"0000000000000000000000001000000000000000000000000000000000000000",
		INIT_27 => X"0000000000000000000000000000000000100000200003000000000002000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2D => X"0000000000000000000000000000000000000000009000900000000000000000",
		INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2F => X"0000000099999999000000000000000000000000000000000000000000000000",
		INIT_30 => X"0000000000000000000000000000000000000000000000000000000000999900",
		INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"5555555500000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"0000515551154000001150155155550000114555514515000000000000000000",
		INIT_39 => X"0000000000000000000000000000000000000015455000000001555451545400",
		INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"550005000000055500555505555500000000000000000000ffc00c00c03cc300"
	)
	port map (
		CLKA => clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(7 downto 7),
		DOA => cpu_D_out(7 downto 7),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(7 downto 7),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

end Behavioral;
